/*
ALUctr[3]	ALUctr[2:0]}	ALU操作

0	        0	            选择加法器输出，做加法
1	        0	            选择加法器输出，做减法
×	        1	            选择移位器输出，左移
0	        10	            做减法，选择带符号小于置位结果输出, Less按带符号结果设置
1	        10	            做减法，选择无符号小于置位结果输出, Less按无符号结果设置
×	        11	            选择ALU输入B的结果直接输出
×	        100	            选择异或输出
0	        101	            选择移位器输出，逻辑右移
1	        101	            选择移位器输出，算术右移
×	        110	            选择逻辑或输出
×	        111	            选择逻辑与输出
*/


module ALU(
        input [31:0] A,
        input [31:0] B,
        input [3:0] ctr,
        output [31:0] out
    );

    assign out = A + B;

endmodule
